library ieee;
	use ieee.std_logic_1164.all;
	use ieee.numeric_std.all;


package filter_pkg is

	type coefficient_array is array(natural range <>) of real;
	type natural_array     is array(natural range <>) of natural;

end package;

package body filter_pkg is

end package body;
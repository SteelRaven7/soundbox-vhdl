----------------------------------
-- testbench type 3 for         --
-- multiplier/accumulator (MAC) --
-- for generic vector           --
----------------------------------

LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
USE ieee.numeric_std.ALL;

ENTITY decimator_tb IS
   
   PORT(y:OUT STD_LOGIC_VECTOR(15 DOWNTO 0)  );
END decimator_tb;

ARCHITECTURE arch_decimator_tb OF
                     decimator_tb IS

   COMPONENT Decimator is
    Port ( input: in std_logic_vector(15 downto 0);
           output: out std_logic_vector(15 downto 0);
           clk :in std_logic;
           reset:in std_logic
            );
           
   END COMPONENT Decimator;

   SIGNAL x_tb_signal:STD_LOGIC_VECTOR(15 DOWNTO 0);
   SIGNAL y_tb_signal:STD_LOGIC_VECTOR(15 DOWNTO 0);
   SIGNAL clk_tb_signal:STD_LOGIC:='0';
   SIGNAL reset_tb_signal:STD_LOGIC;
   
BEGIN
   decimator_comp:
   COMPONENT Decimator
         PORT MAP(clk=>clk_tb_signal,
                  reset=>reset_tb_signal,
                  input=>x_tb_signal,
                  output=>y_tb_signal);
                  
   
    y <= y_tb_signal;

   reset_tb_signal<='0',
                    '1' AFTER 15 ns,
                    '0' AFTER 25 ns;

   
   x_tb_signal<="0000000000000000",  -- 0
                "0001000100010000" AFTER 20 ns, -- 0,5=64
                "0010001000100000" AFTER 40 ns, -- -0,25=-32=224
                "0011001100110000" AFTER 60 ns, -- 0,375=48
                "0100010001000000" AFTER 80 ns, -- -0,75=-96=160
                "0101010101010000" AFTER 100 ns, -- -0,25=-32=224
                "0110011001100000" AFTER 120 ns, -- 0,375=48
                "0111011101110000" AFTER 140 ns, -- -0,75=-96=160
                "1000100010000000" AFTER 160 ns,
                "1001100110010000" AFTER 180 ns,
                "1010101010100000" AFTER 200 ns,
                "1011101110110000" AFTER 220 ns,
                "1100110011000000" AFTER 240 ns,
                "1101110111010000" AFTER 260 ns,
                "1110111011100000" AFTER 280 ns,
                "1111111111110000" AFTER 300 ns,
                "0000000000000000" AFTER 320 ns,
                "0001000100010000" AFTER 340 ns, -- 0,5=64
                "0010001000100000" AFTER 360 ns, -- -0,25=-32=224
                "0011001100110000" AFTER 380 ns, -- 0,375=48
                "0100010001000000" AFTER 400 ns, -- -0,75=-96=160
                "0101010101010000" AFTER 420 ns, -- -0,25=-32=224
                "0110011001100000" AFTER 440 ns, -- 0,375=48
                "0111011101110000" AFTER 460 ns, -- -0,75=-96=160
                "1000100010000000" AFTER 480 ns,
                "1001100110010000" AFTER 500 ns,
                "1010101010100000" AFTER 520 ns,
                "1011101110110000" AFTER 540 ns,
                "1100110011000000" AFTER 560 ns,
                "1101110111010000" AFTER 580 ns,
                "1110111011100000" AFTER 600 ns,
                "1111111111110000" AFTER 620 ns,
                "0000000000000000" AFTER 640 ns,
                "0001000100010000" AFTER 660 ns, -- 0,5=64
                "0010001000100000" AFTER 680 ns, -- -0,25=-32=224
                "0011001100110000" AFTER 700 ns, -- 0,375=48
                "0100010001000000" AFTER 720 ns, -- -0,75=-96=160
                "0101010101010000" AFTER 740 ns, -- -0,25=-32=224
                "0110011001100000" AFTER 760 ns, -- 0,375=48
                "0111011101110000" AFTER 780 ns, -- -0,75=-96=160
                "1000100010000000" AFTER 800 ns,
                "1001100110010000" AFTER 820 ns,
                "1010101010100000" AFTER 840 ns,
                "1011101110110000" AFTER 860 ns,
                "1100110011000000" AFTER 880 ns,
                "1101110111010000" AFTER 900 ns,
                "1110111011100000" AFTER 920 ns, 
                "1111111111110000" AFTER 940 ns,
                "0000000000000000" AFTER 960 ns,
                "0001000100010000" AFTER 980 ns, -- 0,5=64
                "0010001000100000" AFTER 1000 ns, -- -0,25=-32=224
                "0011001100110000" AFTER 1020 ns, -- 0,375=48
                "0100010001000000" AFTER 1040 ns, -- -0,75=-96=160
                "0101010101010000" AFTER 1060 ns, -- -0,25=-32=224
                "0110011001100000" AFTER 1080 ns, -- 0,375=48
                "0111011101110000" AFTER 1100 ns, -- -0,75=-96=160
                "1000100010000000" AFTER 1120 ns,
                "1001100110010000" AFTER 1140 ns,
                "1010101010100000" AFTER 1160 ns,
                "1011101110110000" AFTER 1180 ns,
                "1100110011000000" AFTER 1200 ns,
                "1101110111010000" AFTER 1220 ns,
                "1110111011100000" AFTER 1240 ns,
                "1111111111110000" AFTER 1260 ns,
                "0000000000000000" AFTER 1280 ns,  -- 0
                "0001000100010000" AFTER 1300 ns, -- 0,5=64
                "0010001000100000" AFTER 1320 ns, -- -0,25=-32=224
                "0011001100110000" AFTER 1340 ns, -- 0,375=48
                "0100010001000000" AFTER 1360 ns, -- -0,75=-96=160
                "0101010101010000" AFTER 1380 ns, -- -0,25=-32=224
                "0110011001100000" AFTER 1400 ns, -- 0,375=48
                "0111011101110000" AFTER 1420 ns, -- -0,75=-96=160
                "1000100010000000" AFTER 1440 ns,
                "1001100110010000" AFTER 1460 ns,
                "1010101010100000" AFTER 1480 ns,
                "1011101110110000" AFTER 1500 ns,
                "1100110011000000" AFTER 1520 ns,
                "1101110111010000" AFTER 1540 ns,
                "1110111011100000" AFTER 1560 ns,
                "1111111111110000" AFTER 1580 ns,
                "0000000000000000" AFTER 1600 ns,
                "0001000100010000" AFTER 1620 ns, -- 0,5=64
                "0010001000100000" AFTER 1640 ns, -- -0,25=-32=224
                "0011001100110000" AFTER 1660 ns, -- 0,375=48
                "0100010001000000" AFTER 1680 ns, -- -0,75=-96=160
                "0101010101010000" AFTER 1700 ns, -- -0,25=-32=224
                "0110011001100000" AFTER 1720 ns, -- 0,375=48
                "0111011101110000" AFTER 1740 ns, -- -0,75=-96=160
                "1000100010000000" AFTER 1760 ns,
                "1001100110010000" AFTER 1780 ns,
                "1010101010100000" AFTER 1800 ns,
                "1011101110110000" AFTER 1820 ns,
                "1100110011000000" AFTER 1840 ns,
                "1101110111010000" AFTER 1860 ns,
                "1110111011100000" AFTER 1880 ns,
                "1111111111110000" AFTER 1900 ns,
                "0000000000000000" AFTER 1920 ns,
                "0001000100010000" AFTER 1940 ns, -- 0,5=64
                "0010001000100000" AFTER 1960 ns, -- -0,25=-32=224
                "0011001100110000" AFTER 1980 ns, -- 0,375=48
                "0100010001000000" AFTER 2000 ns, -- -0,75=-96=160
                "0101010101010000" AFTER 2020 ns, -- -0,25=-32=224
                "0110011001100000" AFTER 2040 ns, -- 0,375=48
                "0111011101110000" AFTER 2060 ns, -- -0,75=-96=160
                "1000100010000000" AFTER 2080 ns,
                "1001100110010000" AFTER 2100 ns,
                "1010101010100000" AFTER 2120 ns,
                "1011101110110000" AFTER 2140 ns,
                "1100110011000000" AFTER 2160 ns,
                "1101110111010000" AFTER 2180 ns,
                "1110111011100000" AFTER 2200 ns, 
                "1111111111110000" AFTER 2220 ns,
                "0000000000000000" AFTER 2240 ns,
                "0001000100010000" AFTER 2260 ns, -- 0,5=64
                "0010001000100000" AFTER 2280 ns, -- -0,25=-32=224
                "0011001100110000" AFTER 2300 ns, -- 0,375=48
                "0100010001000000" AFTER 2320 ns, -- -0,75=-96=160
                "0101010101010000" AFTER 2340 ns, -- -0,25=-32=224
                "0110011001100000" AFTER 2360 ns, -- 0,375=48
                "0111011101110000" AFTER 2380 ns, -- -0,75=-96=160
                "1000100010000000" AFTER 2400 ns,
                "1001100110010000" AFTER 2420 ns,
                "1010101010100000" AFTER 2440 ns,
                "1011101110110000" AFTER 2460 ns,
                "1100110011000000" AFTER 2480 ns,
                "1101110111010000" AFTER 2500 ns,
                "1110111011100000" AFTER 2520 ns,
                "1111111111110000" AFTER 2540 ns,
                "0000000000000000" AFTER 2560 ns,  -- 0
                "0001000100010000" AFTER 2580 ns, -- 0,5=64
                "0010001000100000" AFTER 2600 ns, -- -0,25=-32=224
                "0011001100110000" AFTER 2620 ns, -- 0,375=48
                "0100010001000000" AFTER 2640 ns, -- -0,75=-96=160
                "0101010101010000" AFTER 2660 ns, -- -0,25=-32=224
                "0110011001100000" AFTER 2680 ns, -- 0,375=48
                "0111011101110000" AFTER 2700 ns, -- -0,75=-96=160
                "1000100010000000" AFTER 2720 ns,
                "1001100110010000" AFTER 2740 ns,
                "1010101010100000" AFTER 2760 ns,
                "1011101110110000" AFTER 2780 ns,
                "1100110011000000" AFTER 2800 ns,
                "1101110111010000" AFTER 2820 ns,
                "1110111011100000" AFTER 2840 ns,
                "1111111111110000" AFTER 2860 ns,
                "0000000000000000" AFTER 2880 ns,
                "0001000100010000" AFTER 2900 ns, -- 0,5=64
                "0010001000100000" AFTER 2920 ns, -- -0,25=-32=224
                "0011001100110000" AFTER 2940 ns, -- 0,375=48
                "0100010001000000" AFTER 2960 ns, -- -0,75=-96=160
                "0101010101010000" AFTER 2980 ns, -- -0,25=-32=224
                "0110011001100000" AFTER 3000 ns, -- 0,375=48
                "0111011101110000" AFTER 3020 ns, -- -0,75=-96=160
                "1000100010000000" AFTER 3040 ns,
                "1001100110010000" AFTER 3060 ns,
                "1010101010100000" AFTER 3080 ns,
                "1011101110110000" AFTER 3100 ns,
                "1100110011000000" AFTER 3120 ns,
                "1101110111010000" AFTER 3140 ns,
                "1110111011100000" AFTER 3160 ns,
                "1111111111110000" AFTER 3180 ns,
                "0000000000000000" AFTER 3200 ns,
                "0001000100010000" AFTER 3220 ns, -- 0,5=64
                "0010001000100000" AFTER 3240 ns, -- -0,25=-32=224
                "0011001100110000" AFTER 3260 ns, -- 0,375=48
                "0100010001000000" AFTER 3280 ns, -- -0,75=-96=160
                "0101010101010000" AFTER 3300 ns, -- -0,25=-32=224
                "0110011001100000" AFTER 3320 ns, -- 0,375=48
                "0111011101110000" AFTER 3340 ns, -- -0,75=-96=160
                "1000100010000000" AFTER 3360 ns,
                "1001100110010000" AFTER 3380 ns,
                "1010101010100000" AFTER 3400 ns,
                "1011101110110000" AFTER 3420 ns,
                "1100110011000000" AFTER 3440 ns,
                "1101110111010000" AFTER 3460 ns,
                "1110111011100000" AFTER 3480 ns, 
                "1111111111110000" AFTER 3500 ns,
                "0000000000000000" AFTER 3520 ns,
                "0001000100010000" AFTER 3540 ns, -- 0,5=64
                "0010001000100000" AFTER 3560 ns, -- -0,25=-32=224
                "0011001100110000" AFTER 3580 ns, -- 0,375=48
                "0100010001000000" AFTER 3600 ns, -- -0,75=-96=160
                "0101010101010000" AFTER 3620 ns, -- -0,25=-32=224
                "0110011001100000" AFTER 3640 ns, -- 0,375=48
                "0111011101110000" AFTER 3660 ns, -- -0,75=-96=160
                "1000100010000000" AFTER 3680 ns,
                "1001100110010000" AFTER 3700 ns,
                "1010101010100000" AFTER 3720 ns,
                "1011101110110000" AFTER 3740 ns,
                "1100110011000000" AFTER 3760 ns,
                "1101110111010000" AFTER 3780 ns,
                "1110111011100000" AFTER 3800 ns,
                "1111111111110000" AFTER 3820 ns,
                "0000000000000000" AFTER 3840 ns,  -- 0
                "0001000100010000" AFTER 3860 ns, -- 0,5=64
                "0010001000100000" AFTER 3880 ns, -- -0,25=-32=224
                "0011001100110000" AFTER 3900 ns, -- 0,375=48
                "0100010001000000" AFTER 3920 ns, -- -0,75=-96=160
                "0101010101010000" AFTER 3940 ns, -- -0,25=-32=224
                "0110011001100000" AFTER 3960 ns, -- 0,375=48
                "0111011101110000" AFTER 3980 ns, -- -0,75=-96=160
                "1000100010000000" AFTER 4000 ns,
                "1001100110010000" AFTER 4020 ns,
                "1010101010100000" AFTER 4040 ns,
                "1011101110110000" AFTER 4060 ns,
                "1100110011000000" AFTER 4080 ns,
                "1101110111010000" AFTER 4100 ns,
                "1110111011100000" AFTER 4120 ns,
                "1111111111110000" AFTER 4140 ns,
                "0000000000000000" AFTER 4160 ns,
                "0001000100010000" AFTER 4180 ns, -- 0,5=64
                "0010001000100000" AFTER 4200 ns, -- -0,25=-32=224
                "0011001100110000" AFTER 4220 ns, -- 0,375=48
                "0100010001000000" AFTER 4240 ns, -- -0,75=-96=160
                "0101010101010000" AFTER 4260 ns, -- -0,25=-32=224
                "0110011001100000" AFTER 4280 ns, -- 0,375=48
                "0111011101110000" AFTER 4300 ns, -- -0,75=-96=160
                "1000100010000000" AFTER 4320 ns,
                "1001100110010000" AFTER 4340 ns,
                "1010101010100000" AFTER 4360 ns,
                "1011101110110000" AFTER 4380 ns,
                "1100110011000000" AFTER 4400 ns,
                "1101110111010000" AFTER 4420 ns,
                "1110111011100000" AFTER 4440 ns,
                "1111111111110000" AFTER 4460 ns,
                "0000000000000000" AFTER 4480 ns,
                "0001000100010000" AFTER 4500 ns, -- 0,5=64
                "0010001000100000" AFTER 4520 ns, -- -0,25=-32=224
                "0011001100110000" AFTER 4540 ns, -- 0,375=48
                "0100010001000000" AFTER 4560 ns, -- -0,75=-96=160
                "0101010101010000" AFTER 4580 ns, -- -0,25=-32=224
                "0110011001100000" AFTER 4600 ns, -- 0,375=48
                "0111011101110000" AFTER 4620 ns, -- -0,75=-96=160
                "1000100010000000" AFTER 4640 ns,
                "1001100110010000" AFTER 4660 ns,
                "1010101010100000" AFTER 4680 ns,
                "1011101110110000" AFTER 4700 ns,
                "1100110011000000" AFTER 4720 ns,
                "1101110111010000" AFTER 4740 ns,
                "1110111011100000" AFTER 4760 ns, 
                "1111111111110000" AFTER 4780 ns,
                "0000000000000000" AFTER 4800 ns,
                "0001000100010000" AFTER 4820 ns, -- 0,5=64
                "0010001000100000" AFTER 4840 ns, -- -0,25=-32=224
                "0011001100110000" AFTER 4860 ns, -- 0,375=48
                "0100010001000000" AFTER 4880 ns, -- -0,75=-96=160
                "0101010101010000" AFTER 4900 ns, -- -0,25=-32=224
                "0110011001100000" AFTER 4920 ns, -- 0,375=48
                "0111011101110000" AFTER 4940 ns, -- -0,75=-96=160
                "1000100010000000" AFTER 4960 ns,
                "1001100110010000" AFTER 4980 ns,
                "1010101010100000" AFTER 5000 ns,
                "1011101110110000" AFTER 5020 ns,
                "1100110011000000" AFTER 5040 ns,
                "1101110111010000" AFTER 5060 ns,
                "1110111011100000" AFTER 5080 ns,
                "1111111111110000" AFTER 5100 ns;
   clock_proc: process
   begin
      WAIT FOR 10 ns;
      clk_tb_signal<=NOT(clk_tb_signal);
   end process clock_proc ;

  END arch_decimator_tb;